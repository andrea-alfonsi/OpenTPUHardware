`include "rtl/core/control/instruction_decoder.sv"

module instruction_decoder_tb;
  logic clk = 0;

  instruction_decoder id( .* );  
endmodule
