module dut(input a, input b, output o);
  assign o = a ^ b;
endmodule