// todo
`include "rtl/core/systolic_arrays/roundabout_systolic_array.sv"

module roundabout_systolic_array_tb;

endmodule